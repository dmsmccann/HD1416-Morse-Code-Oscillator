.title KiCad schematic
.include "Pot.lib"
.include "Pot2.lib"
.include "standard.bjt"
.include "standard.dio"
V1 +9 GND dc 9
D1 GND Net-_C1-Pad1_ D1N4005
C1 Net-_C1-Pad1_ GND .01u
Q2 /astable2 /node6 GND MPSA20
C4 /astable2 Net-_C4-Pad2_ .1u
R5 +9 /astable2 5.6k
R4 Net-_R3-Pad2_ /node6 68k
R6 Net-_C5-Pad2_ GND 2.2k
XR8 Net-_C4-Pad2_ Net-_C5-Pad1_ GND pot_lin
RJ1 Net-_H3-Pad1_ Net-_C5-Pad1_ 1
R9 GND Net-_H3-Pad1_ 8200
C5 Net-_C5-Pad1_ Net-_C5-Pad2_ .2u
RLS1 +9 /speaker 50
R7 +9 Net-_C5-Pad2_ 33k
Q3 /speaker Net-_C5-Pad2_ GND BC547A
C2 /astable2 /node5 .005u
R2 +9 /node5 220k
C3 /astable1 /node6 .01u
Q1 /astable1 /node5 GND MPSA20
R1 +9 /astable1 10k
XR3 +9 Net-_R3-Pad2_ GND pot_lin2
.param Rt=25k set=0.5 Rt2=500k set2=0.5
.tran 1u 50m 0
.end
